module part1 (
  input [31:0] numbers[4095:0]; // assuming a maximum of 4096 numbers
  output [31:0] out;
);
  
endmodule


